`timescale 1ns/1ps
module MUX81(
    output wire [7:0]o,
    input wire [7:0][7:0]i,
    input wire [2:0]s
);

    wire [7:0][7:0]mins;
    wire [2:0] ns;
    not n0(ns[0],s[0]);
    not n1(ns[1],s[1]);
    not n2(ns[2],s[2]);
    wire [7:0] s1;
    and a0(s1[0],ns[0],ns[1],ns[2]);
    and a1(s1[1],s[0],ns[1],ns[2]);
    and a2(s1[2],ns[0],s[1],ns[2]);
    and a3(s1[3],s[0],s[1],ns[2]);
    and a4(s1[4],ns[0],ns[1],s[2]);
    and a5(s1[5],s[0],ns[1],s[2]);
    and a6(s1[6],ns[0],s[1],s[2]);
    and a7(s1[7],s[0],s[1],s[2]);

and aa10(mins[0][0],s1[0],i[0][0]);
and aa11(mins[0][1],s1[0],i[0][1]);
and aa12(mins[0][2],s1[0],i[0][2]);
and aa13(mins[0][3],s1[0],i[0][3]);
and aa14(mins[0][4],s1[0],i[0][4]);
and aa15(mins[0][5],s1[0],i[0][5]);
and aa16(mins[0][6],s1[0],i[0][6]);
and aa17(mins[0][7],s1[0],i[0][7]);

and aa20(mins[1][0],s1[1],i[1][0]);
and aa21(mins[1][1],s1[1],i[1][1]);
and aa22(mins[1][2],s1[1],i[1][2]);
and aa23(mins[1][3],s1[1],i[1][3]);
and aa24(mins[1][4],s1[1],i[1][4]);
and aa25(mins[1][5],s1[1],i[1][5]);
and aa26(mins[1][6],s1[1],i[1][6]);
and aa27(mins[1][7],s1[1],i[1][7]);

and aa30(mins[2][0],s1[2],i[2][0]);
and aa31(mins[2][1],s1[2],i[2][1]);
and aa32(mins[2][2],s1[2],i[2][2]);
and aa33(mins[2][3],s1[2],i[2][3]);
and aa34(mins[2][4],s1[2],i[2][4]);
and aa35(mins[2][5],s1[2],i[2][5]);
and aa36(mins[2][6],s1[2],i[2][6]);
and aa37(mins[2][7],s1[2],i[2][7]);

and aa40(mins[3][0],s1[3],i[3][0]);
and aa41(mins[3][1],s1[3],i[3][1]);
and aa42(mins[3][2],s1[3],i[3][2]);
and aa43(mins[3][3],s1[3],i[3][3]);
and aa44(mins[3][4],s1[3],i[3][4]);
and aa45(mins[3][5],s1[3],i[3][5]);
and aa46(mins[3][6],s1[3],i[3][6]);
and aa47(mins[3][7],s1[3],i[3][7]);

and aa50(mins[4][0],s1[4],i[4][0]);
and aa51(mins[4][1],s1[4],i[4][1]);
and aa52(mins[4][2],s1[4],i[4][2]);
and aa53(mins[4][3],s1[4],i[4][3]);
and aa54(mins[4][4],s1[4],i[4][4]);
and aa55(mins[4][5],s1[4],i[4][5]);
and aa56(mins[4][6],s1[4],i[4][6]);
and aa57(mins[4][7],s1[4],i[4][7]);

and aa60(mins[5][0],s1[5],i[5][0]);
and aa61(mins[5][1],s1[5],i[5][1]);
and aa62(mins[5][2],s1[5],i[5][2]);
and aa63(mins[5][3],s1[5],i[5][3]);
and aa64(mins[5][4],s1[5],i[5][4]);
and aa65(mins[5][5],s1[5],i[5][5]);
and aa66(mins[5][6],s1[5],i[5][6]);
and aa67(mins[5][7],s1[5],i[5][7]);

and aa70(mins[6][0],s1[6],i[6][0]);
and aa71(mins[6][1],s1[6],i[6][1]);
and aa72(mins[6][2],s1[6],i[6][2]);
and aa73(mins[6][3],s1[6],i[6][3]);
and aa74(mins[6][4],s1[6],i[6][4]);
and aa75(mins[6][5],s1[6],i[6][5]);
and aa76(mins[6][6],s1[6],i[6][6]);
and aa77(mins[6][7],s1[6],i[6][7]);

and aa80(mins[7][0],s1[7],i[7][0]);
and aa81(mins[7][1],s1[7],i[7][1]);
and aa82(mins[7][2],s1[7],i[7][2]);
and aa83(mins[7][3],s1[7],i[7][3]);
and aa84(mins[7][4],s1[7],i[7][4]);
and aa85(mins[7][5],s1[7],i[7][5]);
and aa86(mins[7][6],s1[7],i[7][6]);
and aa87(mins[7][7],s1[7],i[7][7]);

or op0(o[0],mins[0][0],mins[1][0],mins[2][0],mins[3][0],mins[4][0],mins[5][0],mins[6][0],mins[7][0]);
or op1(o[1],mins[0][1],mins[1][1],mins[2][1],mins[3][1],mins[4][1],mins[5][1],mins[6][1],mins[7][1]);
or op2(o[2],mins[0][2],mins[1][2],mins[2][2],mins[3][2],mins[4][2],mins[5][2],mins[6][2],mins[7][2]);
or op3(o[3],mins[0][3],mins[1][3],mins[2][3],mins[3][3],mins[4][3],mins[5][3],mins[6][3],mins[7][3]);
or op4(o[4],mins[0][4],mins[1][4],mins[2][4],mins[3][4],mins[4][4],mins[5][4],mins[6][4],mins[7][4]);
or op5(o[5],mins[0][5],mins[1][5],mins[2][5],mins[3][5],mins[4][5],mins[5][5],mins[6][5],mins[7][5]);
or op6(o[6],mins[0][6],mins[1][6],mins[2][6],mins[3][6],mins[4][6],mins[5][6],mins[6][6],mins[7][6]);
or op7(o[7],mins[0][7],mins[1][7],mins[2][7],mins[3][7],mins[4][7],mins[5][7],mins[6][7],mins[7][7]);

endmodule